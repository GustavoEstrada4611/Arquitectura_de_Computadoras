//1. Definicion de modulo y sus entradas y salidas
module _and (input A, input B, output C);
//2. Declarar señales/elementos internos
//NA
//3. Comportamiento del modulo
	//(Asignaciones, Instancias, Conexiones)
assign C=A&B;



endmodule

//Repositorio GitHub: https://github.com/GustavoEstrada4611/Arquitectura_de_Computadoras